library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.math_real.all;

library work;
use work.DFTTypes.all;

package DFTSinusoidLUT is
    
    type sinusoid_LUT_array is   array (2*K_LENGTH-1 downto 0) of signed_fxp_sinusoid;
    
    -- format:
    -- 0: cos(-2*pi*k0/#samples)
    -- 1: sin(-2*pi*k0/#samples)
    -- 2: cos(-2*pi*k1/#samples)
    -- 3: sin(-2*pi*k1/#samples)
    -- ...

    constant K_SINUSOID_LUT   : sinusoid_LUT_array :=
        (
            to_signed(32767, signed_fxp_sinusoid'length),
            to_signed(0, signed_fxp_sinusoid'length),
            to_signed(32765, signed_fxp_sinusoid'length),
            to_signed(-402, signed_fxp_sinusoid'length),
            to_signed(32758, signed_fxp_sinusoid'length),
            to_signed(-804, signed_fxp_sinusoid'length),
            to_signed(32745, signed_fxp_sinusoid'length),
            to_signed(-1206, signed_fxp_sinusoid'length),
            to_signed(32728, signed_fxp_sinusoid'length),
            to_signed(-1607, signed_fxp_sinusoid'length),
            to_signed(32706, signed_fxp_sinusoid'length),
            to_signed(-2009, signed_fxp_sinusoid'length),
            to_signed(32679, signed_fxp_sinusoid'length),
            to_signed(-2410, signed_fxp_sinusoid'length),
            to_signed(32647, signed_fxp_sinusoid'length),
            to_signed(-2811, signed_fxp_sinusoid'length),
            to_signed(32610, signed_fxp_sinusoid'length),
            to_signed(-3211, signed_fxp_sinusoid'length),
            to_signed(32568, signed_fxp_sinusoid'length),
            to_signed(-3611, signed_fxp_sinusoid'length),
            to_signed(32521, signed_fxp_sinusoid'length),
            to_signed(-4011, signed_fxp_sinusoid'length),
            to_signed(32469, signed_fxp_sinusoid'length),
            to_signed(-4409, signed_fxp_sinusoid'length),
            to_signed(32413, signed_fxp_sinusoid'length),
            to_signed(-4808, signed_fxp_sinusoid'length),
            to_signed(32351, signed_fxp_sinusoid'length),
            to_signed(-5205, signed_fxp_sinusoid'length),
            to_signed(32285, signed_fxp_sinusoid'length),
            to_signed(-5602, signed_fxp_sinusoid'length),
            to_signed(32214, signed_fxp_sinusoid'length),
            to_signed(-5997, signed_fxp_sinusoid'length),
            to_signed(32138, signed_fxp_sinusoid'length),
            to_signed(-6392, signed_fxp_sinusoid'length),
            to_signed(32057, signed_fxp_sinusoid'length),
            to_signed(-6786, signed_fxp_sinusoid'length),
            to_signed(31971, signed_fxp_sinusoid'length),
            to_signed(-7179, signed_fxp_sinusoid'length),
            to_signed(31881, signed_fxp_sinusoid'length),
            to_signed(-7571, signed_fxp_sinusoid'length),
            to_signed(31785, signed_fxp_sinusoid'length),
            to_signed(-7961, signed_fxp_sinusoid'length),
            to_signed(31685, signed_fxp_sinusoid'length),
            to_signed(-8351, signed_fxp_sinusoid'length),
            to_signed(31581, signed_fxp_sinusoid'length),
            to_signed(-8739, signed_fxp_sinusoid'length),
            to_signed(31471, signed_fxp_sinusoid'length),
            to_signed(-9126, signed_fxp_sinusoid'length),
            to_signed(31357, signed_fxp_sinusoid'length),
            to_signed(-9512, signed_fxp_sinusoid'length),
            to_signed(31237, signed_fxp_sinusoid'length),
            to_signed(-9896, signed_fxp_sinusoid'length),
            to_signed(31114, signed_fxp_sinusoid'length),
            to_signed(-10278, signed_fxp_sinusoid'length),
            to_signed(30985, signed_fxp_sinusoid'length),
            to_signed(-10659, signed_fxp_sinusoid'length),
            to_signed(30852, signed_fxp_sinusoid'length),
            to_signed(-11039, signed_fxp_sinusoid'length),
            to_signed(30714, signed_fxp_sinusoid'length),
            to_signed(-11416, signed_fxp_sinusoid'length),
            to_signed(30572, signed_fxp_sinusoid'length),
            to_signed(-11793, signed_fxp_sinusoid'length),
            to_signed(30425, signed_fxp_sinusoid'length),
            to_signed(-12167, signed_fxp_sinusoid'length),
            to_signed(30273, signed_fxp_sinusoid'length),
            to_signed(-12539, signed_fxp_sinusoid'length),
            to_signed(30117, signed_fxp_sinusoid'length),
            to_signed(-12910, signed_fxp_sinusoid'length),
            to_signed(29956, signed_fxp_sinusoid'length),
            to_signed(-13278, signed_fxp_sinusoid'length),
            to_signed(29791, signed_fxp_sinusoid'length),
            to_signed(-13645, signed_fxp_sinusoid'length),
            to_signed(29621, signed_fxp_sinusoid'length),
            to_signed(-14010, signed_fxp_sinusoid'length),
            to_signed(29447, signed_fxp_sinusoid'length),
            to_signed(-14372, signed_fxp_sinusoid'length),
            to_signed(29269, signed_fxp_sinusoid'length),
            to_signed(-14732, signed_fxp_sinusoid'length),
            to_signed(29086, signed_fxp_sinusoid'length),
            to_signed(-15090, signed_fxp_sinusoid'length),
            to_signed(28898, signed_fxp_sinusoid'length),
            to_signed(-15446, signed_fxp_sinusoid'length),
            to_signed(28707, signed_fxp_sinusoid'length),
            to_signed(-15800, signed_fxp_sinusoid'length),
            to_signed(28511, signed_fxp_sinusoid'length),
            to_signed(-16151, signed_fxp_sinusoid'length),
            to_signed(28310, signed_fxp_sinusoid'length),
            to_signed(-16499, signed_fxp_sinusoid'length),
            to_signed(28106, signed_fxp_sinusoid'length),
            to_signed(-16846, signed_fxp_sinusoid'length),
            to_signed(27897, signed_fxp_sinusoid'length),
            to_signed(-17189, signed_fxp_sinusoid'length),
            to_signed(27684, signed_fxp_sinusoid'length),
            to_signed(-17530, signed_fxp_sinusoid'length),
            to_signed(27466, signed_fxp_sinusoid'length),
            to_signed(-17869, signed_fxp_sinusoid'length),
            to_signed(27245, signed_fxp_sinusoid'length),
            to_signed(-18204, signed_fxp_sinusoid'length),
            to_signed(27020, signed_fxp_sinusoid'length),
            to_signed(-18537, signed_fxp_sinusoid'length),
            to_signed(26790, signed_fxp_sinusoid'length),
            to_signed(-18868, signed_fxp_sinusoid'length),
            to_signed(26557, signed_fxp_sinusoid'length),
            to_signed(-19195, signed_fxp_sinusoid'length),
            to_signed(26319, signed_fxp_sinusoid'length),
            to_signed(-19519, signed_fxp_sinusoid'length),
            to_signed(26077, signed_fxp_sinusoid'length),
            to_signed(-19841, signed_fxp_sinusoid'length),
            to_signed(25832, signed_fxp_sinusoid'length),
            to_signed(-20159, signed_fxp_sinusoid'length),
            to_signed(25583, signed_fxp_sinusoid'length),
            to_signed(-20475, signed_fxp_sinusoid'length),
            to_signed(25330, signed_fxp_sinusoid'length),
            to_signed(-20787, signed_fxp_sinusoid'length),
            to_signed(25073, signed_fxp_sinusoid'length),
            to_signed(-21097, signed_fxp_sinusoid'length),
            to_signed(24812, signed_fxp_sinusoid'length),
            to_signed(-21403, signed_fxp_sinusoid'length),
            to_signed(24547, signed_fxp_sinusoid'length),
            to_signed(-21706, signed_fxp_sinusoid'length),
            to_signed(24279, signed_fxp_sinusoid'length),
            to_signed(-22005, signed_fxp_sinusoid'length),
            to_signed(24007, signed_fxp_sinusoid'length),
            to_signed(-22301, signed_fxp_sinusoid'length),
            to_signed(23732, signed_fxp_sinusoid'length),
            to_signed(-22594, signed_fxp_sinusoid'length),
            to_signed(23453, signed_fxp_sinusoid'length),
            to_signed(-22884, signed_fxp_sinusoid'length),
            to_signed(23170, signed_fxp_sinusoid'length),
            to_signed(-23170, signed_fxp_sinusoid'length),
            to_signed(22884, signed_fxp_sinusoid'length),
            to_signed(-23453, signed_fxp_sinusoid'length),
            to_signed(22594, signed_fxp_sinusoid'length),
            to_signed(-23732, signed_fxp_sinusoid'length),
            to_signed(22301, signed_fxp_sinusoid'length),
            to_signed(-24007, signed_fxp_sinusoid'length),
            to_signed(22005, signed_fxp_sinusoid'length),
            to_signed(-24279, signed_fxp_sinusoid'length),
            to_signed(21706, signed_fxp_sinusoid'length),
            to_signed(-24547, signed_fxp_sinusoid'length),
            to_signed(21403, signed_fxp_sinusoid'length),
            to_signed(-24812, signed_fxp_sinusoid'length),
            to_signed(21097, signed_fxp_sinusoid'length),
            to_signed(-25073, signed_fxp_sinusoid'length),
            to_signed(20787, signed_fxp_sinusoid'length),
            to_signed(-25330, signed_fxp_sinusoid'length),
            to_signed(20475, signed_fxp_sinusoid'length),
            to_signed(-25583, signed_fxp_sinusoid'length),
            to_signed(20159, signed_fxp_sinusoid'length),
            to_signed(-25832, signed_fxp_sinusoid'length),
            to_signed(19841, signed_fxp_sinusoid'length),
            to_signed(-26077, signed_fxp_sinusoid'length),
            to_signed(19519, signed_fxp_sinusoid'length),
            to_signed(-26319, signed_fxp_sinusoid'length),
            to_signed(19195, signed_fxp_sinusoid'length),
            to_signed(-26557, signed_fxp_sinusoid'length),
            to_signed(18868, signed_fxp_sinusoid'length),
            to_signed(-26790, signed_fxp_sinusoid'length),
            to_signed(18537, signed_fxp_sinusoid'length),
            to_signed(-27020, signed_fxp_sinusoid'length),
            to_signed(18204, signed_fxp_sinusoid'length),
            to_signed(-27245, signed_fxp_sinusoid'length),
            to_signed(17869, signed_fxp_sinusoid'length),
            to_signed(-27466, signed_fxp_sinusoid'length),
            to_signed(17530, signed_fxp_sinusoid'length),
            to_signed(-27684, signed_fxp_sinusoid'length),
            to_signed(17189, signed_fxp_sinusoid'length),
            to_signed(-27897, signed_fxp_sinusoid'length),
            to_signed(16846, signed_fxp_sinusoid'length),
            to_signed(-28106, signed_fxp_sinusoid'length),
            to_signed(16499, signed_fxp_sinusoid'length),
            to_signed(-28310, signed_fxp_sinusoid'length),
            to_signed(16151, signed_fxp_sinusoid'length),
            to_signed(-28511, signed_fxp_sinusoid'length),
            to_signed(15800, signed_fxp_sinusoid'length),
            to_signed(-28707, signed_fxp_sinusoid'length),
            to_signed(15446, signed_fxp_sinusoid'length),
            to_signed(-28898, signed_fxp_sinusoid'length),
            to_signed(15090, signed_fxp_sinusoid'length),
            to_signed(-29086, signed_fxp_sinusoid'length),
            to_signed(14732, signed_fxp_sinusoid'length),
            to_signed(-29269, signed_fxp_sinusoid'length),
            to_signed(14372, signed_fxp_sinusoid'length),
            to_signed(-29447, signed_fxp_sinusoid'length),
            to_signed(14010, signed_fxp_sinusoid'length),
            to_signed(-29621, signed_fxp_sinusoid'length),
            to_signed(13645, signed_fxp_sinusoid'length),
            to_signed(-29791, signed_fxp_sinusoid'length),
            to_signed(13278, signed_fxp_sinusoid'length),
            to_signed(-29956, signed_fxp_sinusoid'length),
            to_signed(12910, signed_fxp_sinusoid'length),
            to_signed(-30117, signed_fxp_sinusoid'length),
            to_signed(12539, signed_fxp_sinusoid'length),
            to_signed(-30273, signed_fxp_sinusoid'length),
            to_signed(12167, signed_fxp_sinusoid'length),
            to_signed(-30425, signed_fxp_sinusoid'length),
            to_signed(11793, signed_fxp_sinusoid'length),
            to_signed(-30572, signed_fxp_sinusoid'length),
            to_signed(11416, signed_fxp_sinusoid'length),
            to_signed(-30714, signed_fxp_sinusoid'length),
            to_signed(11039, signed_fxp_sinusoid'length),
            to_signed(-30852, signed_fxp_sinusoid'length),
            to_signed(10659, signed_fxp_sinusoid'length),
            to_signed(-30985, signed_fxp_sinusoid'length),
            to_signed(10278, signed_fxp_sinusoid'length),
            to_signed(-31114, signed_fxp_sinusoid'length),
            to_signed(9896, signed_fxp_sinusoid'length),
            to_signed(-31237, signed_fxp_sinusoid'length),
            to_signed(9512, signed_fxp_sinusoid'length),
            to_signed(-31357, signed_fxp_sinusoid'length),
            to_signed(9126, signed_fxp_sinusoid'length),
            to_signed(-31471, signed_fxp_sinusoid'length),
            to_signed(8739, signed_fxp_sinusoid'length),
            to_signed(-31581, signed_fxp_sinusoid'length),
            to_signed(8351, signed_fxp_sinusoid'length),
            to_signed(-31685, signed_fxp_sinusoid'length),
            to_signed(7961, signed_fxp_sinusoid'length),
            to_signed(-31785, signed_fxp_sinusoid'length),
            to_signed(7571, signed_fxp_sinusoid'length),
            to_signed(-31881, signed_fxp_sinusoid'length),
            to_signed(7179, signed_fxp_sinusoid'length),
            to_signed(-31971, signed_fxp_sinusoid'length),
            to_signed(6786, signed_fxp_sinusoid'length),
            to_signed(-32057, signed_fxp_sinusoid'length),
            to_signed(6392, signed_fxp_sinusoid'length),
            to_signed(-32138, signed_fxp_sinusoid'length),
            to_signed(5997, signed_fxp_sinusoid'length),
            to_signed(-32214, signed_fxp_sinusoid'length),
            to_signed(5602, signed_fxp_sinusoid'length),
            to_signed(-32285, signed_fxp_sinusoid'length),
            to_signed(5205, signed_fxp_sinusoid'length),
            to_signed(-32351, signed_fxp_sinusoid'length),
            to_signed(4808, signed_fxp_sinusoid'length),
            to_signed(-32413, signed_fxp_sinusoid'length),
            to_signed(4409, signed_fxp_sinusoid'length),
            to_signed(-32469, signed_fxp_sinusoid'length),
            to_signed(4011, signed_fxp_sinusoid'length),
            to_signed(-32521, signed_fxp_sinusoid'length),
            to_signed(3611, signed_fxp_sinusoid'length),
            to_signed(-32568, signed_fxp_sinusoid'length),
            to_signed(3211, signed_fxp_sinusoid'length),
            to_signed(-32610, signed_fxp_sinusoid'length),
            to_signed(2811, signed_fxp_sinusoid'length),
            to_signed(-32647, signed_fxp_sinusoid'length),
            to_signed(2410, signed_fxp_sinusoid'length),
            to_signed(-32679, signed_fxp_sinusoid'length),
            to_signed(2009, signed_fxp_sinusoid'length),
            to_signed(-32706, signed_fxp_sinusoid'length),
            to_signed(1607, signed_fxp_sinusoid'length),
            to_signed(-32728, signed_fxp_sinusoid'length),
            to_signed(1206, signed_fxp_sinusoid'length),
            to_signed(-32745, signed_fxp_sinusoid'length),
            to_signed(804, signed_fxp_sinusoid'length),
            to_signed(-32758, signed_fxp_sinusoid'length),
            to_signed(402, signed_fxp_sinusoid'length),
            to_signed(-32765, signed_fxp_sinusoid'length),
            to_signed(0, signed_fxp_sinusoid'length),
            to_signed(-32768, signed_fxp_sinusoid'length),
            to_signed(-402, signed_fxp_sinusoid'length),
            to_signed(-32765, signed_fxp_sinusoid'length),
            to_signed(-804, signed_fxp_sinusoid'length),
            to_signed(-32758, signed_fxp_sinusoid'length),
            to_signed(-1206, signed_fxp_sinusoid'length),
            to_signed(-32745, signed_fxp_sinusoid'length),
            to_signed(-1607, signed_fxp_sinusoid'length),
            to_signed(-32728, signed_fxp_sinusoid'length),
            to_signed(-2009, signed_fxp_sinusoid'length),
            to_signed(-32706, signed_fxp_sinusoid'length),
            to_signed(-2410, signed_fxp_sinusoid'length),
            to_signed(-32679, signed_fxp_sinusoid'length),
            to_signed(-2811, signed_fxp_sinusoid'length),
            to_signed(-32647, signed_fxp_sinusoid'length),
            to_signed(-3211, signed_fxp_sinusoid'length),
            to_signed(-32610, signed_fxp_sinusoid'length),
            to_signed(-3611, signed_fxp_sinusoid'length),
            to_signed(-32568, signed_fxp_sinusoid'length),
            to_signed(-4011, signed_fxp_sinusoid'length),
            to_signed(-32521, signed_fxp_sinusoid'length),
            to_signed(-4409, signed_fxp_sinusoid'length),
            to_signed(-32469, signed_fxp_sinusoid'length),
            to_signed(-4808, signed_fxp_sinusoid'length),
            to_signed(-32413, signed_fxp_sinusoid'length),
            to_signed(-5205, signed_fxp_sinusoid'length),
            to_signed(-32351, signed_fxp_sinusoid'length),
            to_signed(-5602, signed_fxp_sinusoid'length),
            to_signed(-32285, signed_fxp_sinusoid'length),
            to_signed(-5997, signed_fxp_sinusoid'length),
            to_signed(-32214, signed_fxp_sinusoid'length),
            to_signed(-6392, signed_fxp_sinusoid'length),
            to_signed(-32138, signed_fxp_sinusoid'length),
            to_signed(-6786, signed_fxp_sinusoid'length),
            to_signed(-32057, signed_fxp_sinusoid'length),
            to_signed(-7179, signed_fxp_sinusoid'length),
            to_signed(-31971, signed_fxp_sinusoid'length),
            to_signed(-7571, signed_fxp_sinusoid'length),
            to_signed(-31881, signed_fxp_sinusoid'length),
            to_signed(-7961, signed_fxp_sinusoid'length),
            to_signed(-31785, signed_fxp_sinusoid'length),
            to_signed(-8351, signed_fxp_sinusoid'length),
            to_signed(-31685, signed_fxp_sinusoid'length),
            to_signed(-8739, signed_fxp_sinusoid'length),
            to_signed(-31581, signed_fxp_sinusoid'length),
            to_signed(-9126, signed_fxp_sinusoid'length),
            to_signed(-31471, signed_fxp_sinusoid'length),
            to_signed(-9512, signed_fxp_sinusoid'length),
            to_signed(-31357, signed_fxp_sinusoid'length),
            to_signed(-9896, signed_fxp_sinusoid'length),
            to_signed(-31237, signed_fxp_sinusoid'length),
            to_signed(-10278, signed_fxp_sinusoid'length),
            to_signed(-31114, signed_fxp_sinusoid'length),
            to_signed(-10659, signed_fxp_sinusoid'length),
            to_signed(-30985, signed_fxp_sinusoid'length),
            to_signed(-11039, signed_fxp_sinusoid'length),
            to_signed(-30852, signed_fxp_sinusoid'length),
            to_signed(-11416, signed_fxp_sinusoid'length),
            to_signed(-30714, signed_fxp_sinusoid'length),
            to_signed(-11793, signed_fxp_sinusoid'length),
            to_signed(-30572, signed_fxp_sinusoid'length),
            to_signed(-12167, signed_fxp_sinusoid'length),
            to_signed(-30425, signed_fxp_sinusoid'length),
            to_signed(-12539, signed_fxp_sinusoid'length),
            to_signed(-30273, signed_fxp_sinusoid'length),
            to_signed(-12910, signed_fxp_sinusoid'length),
            to_signed(-30117, signed_fxp_sinusoid'length),
            to_signed(-13278, signed_fxp_sinusoid'length),
            to_signed(-29956, signed_fxp_sinusoid'length),
            to_signed(-13645, signed_fxp_sinusoid'length),
            to_signed(-29791, signed_fxp_sinusoid'length),
            to_signed(-14010, signed_fxp_sinusoid'length),
            to_signed(-29621, signed_fxp_sinusoid'length),
            to_signed(-14372, signed_fxp_sinusoid'length),
            to_signed(-29447, signed_fxp_sinusoid'length),
            to_signed(-14732, signed_fxp_sinusoid'length),
            to_signed(-29269, signed_fxp_sinusoid'length),
            to_signed(-15090, signed_fxp_sinusoid'length),
            to_signed(-29086, signed_fxp_sinusoid'length),
            to_signed(-15446, signed_fxp_sinusoid'length),
            to_signed(-28898, signed_fxp_sinusoid'length),
            to_signed(-15800, signed_fxp_sinusoid'length),
            to_signed(-28707, signed_fxp_sinusoid'length),
            to_signed(-16151, signed_fxp_sinusoid'length),
            to_signed(-28511, signed_fxp_sinusoid'length),
            to_signed(-16499, signed_fxp_sinusoid'length),
            to_signed(-28310, signed_fxp_sinusoid'length),
            to_signed(-16846, signed_fxp_sinusoid'length),
            to_signed(-28106, signed_fxp_sinusoid'length),
            to_signed(-17189, signed_fxp_sinusoid'length),
            to_signed(-27897, signed_fxp_sinusoid'length),
            to_signed(-17530, signed_fxp_sinusoid'length),
            to_signed(-27684, signed_fxp_sinusoid'length),
            to_signed(-17869, signed_fxp_sinusoid'length),
            to_signed(-27466, signed_fxp_sinusoid'length),
            to_signed(-18204, signed_fxp_sinusoid'length),
            to_signed(-27245, signed_fxp_sinusoid'length),
            to_signed(-18537, signed_fxp_sinusoid'length),
            to_signed(-27020, signed_fxp_sinusoid'length),
            to_signed(-18868, signed_fxp_sinusoid'length),
            to_signed(-26790, signed_fxp_sinusoid'length),
            to_signed(-19195, signed_fxp_sinusoid'length),
            to_signed(-26557, signed_fxp_sinusoid'length),
            to_signed(-19519, signed_fxp_sinusoid'length),
            to_signed(-26319, signed_fxp_sinusoid'length),
            to_signed(-19841, signed_fxp_sinusoid'length),
            to_signed(-26077, signed_fxp_sinusoid'length),
            to_signed(-20159, signed_fxp_sinusoid'length),
            to_signed(-25832, signed_fxp_sinusoid'length),
            to_signed(-20475, signed_fxp_sinusoid'length),
            to_signed(-25583, signed_fxp_sinusoid'length),
            to_signed(-20787, signed_fxp_sinusoid'length),
            to_signed(-25330, signed_fxp_sinusoid'length),
            to_signed(-21097, signed_fxp_sinusoid'length),
            to_signed(-25073, signed_fxp_sinusoid'length),
            to_signed(-21403, signed_fxp_sinusoid'length),
            to_signed(-24812, signed_fxp_sinusoid'length),
            to_signed(-21706, signed_fxp_sinusoid'length),
            to_signed(-24547, signed_fxp_sinusoid'length),
            to_signed(-22005, signed_fxp_sinusoid'length),
            to_signed(-24279, signed_fxp_sinusoid'length),
            to_signed(-22301, signed_fxp_sinusoid'length),
            to_signed(-24007, signed_fxp_sinusoid'length),
            to_signed(-22594, signed_fxp_sinusoid'length),
            to_signed(-23732, signed_fxp_sinusoid'length),
            to_signed(-22884, signed_fxp_sinusoid'length),
            to_signed(-23453, signed_fxp_sinusoid'length),
            to_signed(-23170, signed_fxp_sinusoid'length),
            to_signed(-23170, signed_fxp_sinusoid'length),
            to_signed(-23453, signed_fxp_sinusoid'length),
            to_signed(-22884, signed_fxp_sinusoid'length),
            to_signed(-23732, signed_fxp_sinusoid'length),
            to_signed(-22594, signed_fxp_sinusoid'length),
            to_signed(-24007, signed_fxp_sinusoid'length),
            to_signed(-22301, signed_fxp_sinusoid'length),
            to_signed(-24279, signed_fxp_sinusoid'length),
            to_signed(-22005, signed_fxp_sinusoid'length),
            to_signed(-24547, signed_fxp_sinusoid'length),
            to_signed(-21706, signed_fxp_sinusoid'length),
            to_signed(-24812, signed_fxp_sinusoid'length),
            to_signed(-21403, signed_fxp_sinusoid'length),
            to_signed(-25073, signed_fxp_sinusoid'length),
            to_signed(-21097, signed_fxp_sinusoid'length),
            to_signed(-25330, signed_fxp_sinusoid'length),
            to_signed(-20787, signed_fxp_sinusoid'length),
            to_signed(-25583, signed_fxp_sinusoid'length),
            to_signed(-20475, signed_fxp_sinusoid'length),
            to_signed(-25832, signed_fxp_sinusoid'length),
            to_signed(-20159, signed_fxp_sinusoid'length),
            to_signed(-26077, signed_fxp_sinusoid'length),
            to_signed(-19841, signed_fxp_sinusoid'length),
            to_signed(-26319, signed_fxp_sinusoid'length),
            to_signed(-19519, signed_fxp_sinusoid'length),
            to_signed(-26557, signed_fxp_sinusoid'length),
            to_signed(-19195, signed_fxp_sinusoid'length),
            to_signed(-26790, signed_fxp_sinusoid'length),
            to_signed(-18868, signed_fxp_sinusoid'length),
            to_signed(-27020, signed_fxp_sinusoid'length),
            to_signed(-18537, signed_fxp_sinusoid'length),
            to_signed(-27245, signed_fxp_sinusoid'length),
            to_signed(-18204, signed_fxp_sinusoid'length),
            to_signed(-27466, signed_fxp_sinusoid'length),
            to_signed(-17869, signed_fxp_sinusoid'length),
            to_signed(-27684, signed_fxp_sinusoid'length),
            to_signed(-17530, signed_fxp_sinusoid'length),
            to_signed(-27897, signed_fxp_sinusoid'length),
            to_signed(-17189, signed_fxp_sinusoid'length),
            to_signed(-28106, signed_fxp_sinusoid'length),
            to_signed(-16846, signed_fxp_sinusoid'length),
            to_signed(-28310, signed_fxp_sinusoid'length),
            to_signed(-16499, signed_fxp_sinusoid'length),
            to_signed(-28511, signed_fxp_sinusoid'length),
            to_signed(-16151, signed_fxp_sinusoid'length),
            to_signed(-28707, signed_fxp_sinusoid'length),
            to_signed(-15800, signed_fxp_sinusoid'length),
            to_signed(-28898, signed_fxp_sinusoid'length),
            to_signed(-15446, signed_fxp_sinusoid'length),
            to_signed(-29086, signed_fxp_sinusoid'length),
            to_signed(-15090, signed_fxp_sinusoid'length),
            to_signed(-29269, signed_fxp_sinusoid'length),
            to_signed(-14732, signed_fxp_sinusoid'length),
            to_signed(-29447, signed_fxp_sinusoid'length),
            to_signed(-14372, signed_fxp_sinusoid'length),
            to_signed(-29621, signed_fxp_sinusoid'length),
            to_signed(-14010, signed_fxp_sinusoid'length),
            to_signed(-29791, signed_fxp_sinusoid'length),
            to_signed(-13645, signed_fxp_sinusoid'length),
            to_signed(-29956, signed_fxp_sinusoid'length),
            to_signed(-13278, signed_fxp_sinusoid'length),
            to_signed(-30117, signed_fxp_sinusoid'length),
            to_signed(-12910, signed_fxp_sinusoid'length),
            to_signed(-30273, signed_fxp_sinusoid'length),
            to_signed(-12539, signed_fxp_sinusoid'length),
            to_signed(-30425, signed_fxp_sinusoid'length),
            to_signed(-12167, signed_fxp_sinusoid'length),
            to_signed(-30572, signed_fxp_sinusoid'length),
            to_signed(-11793, signed_fxp_sinusoid'length),
            to_signed(-30714, signed_fxp_sinusoid'length),
            to_signed(-11416, signed_fxp_sinusoid'length),
            to_signed(-30852, signed_fxp_sinusoid'length),
            to_signed(-11039, signed_fxp_sinusoid'length),
            to_signed(-30985, signed_fxp_sinusoid'length),
            to_signed(-10659, signed_fxp_sinusoid'length),
            to_signed(-31114, signed_fxp_sinusoid'length),
            to_signed(-10278, signed_fxp_sinusoid'length),
            to_signed(-31237, signed_fxp_sinusoid'length),
            to_signed(-9896, signed_fxp_sinusoid'length),
            to_signed(-31357, signed_fxp_sinusoid'length),
            to_signed(-9512, signed_fxp_sinusoid'length),
            to_signed(-31471, signed_fxp_sinusoid'length),
            to_signed(-9126, signed_fxp_sinusoid'length),
            to_signed(-31581, signed_fxp_sinusoid'length),
            to_signed(-8739, signed_fxp_sinusoid'length),
            to_signed(-31685, signed_fxp_sinusoid'length),
            to_signed(-8351, signed_fxp_sinusoid'length),
            to_signed(-31785, signed_fxp_sinusoid'length),
            to_signed(-7961, signed_fxp_sinusoid'length),
            to_signed(-31881, signed_fxp_sinusoid'length),
            to_signed(-7571, signed_fxp_sinusoid'length),
            to_signed(-31971, signed_fxp_sinusoid'length),
            to_signed(-7179, signed_fxp_sinusoid'length),
            to_signed(-32057, signed_fxp_sinusoid'length),
            to_signed(-6786, signed_fxp_sinusoid'length),
            to_signed(-32138, signed_fxp_sinusoid'length),
            to_signed(-6392, signed_fxp_sinusoid'length),
            to_signed(-32214, signed_fxp_sinusoid'length),
            to_signed(-5997, signed_fxp_sinusoid'length),
            to_signed(-32285, signed_fxp_sinusoid'length),
            to_signed(-5602, signed_fxp_sinusoid'length),
            to_signed(-32351, signed_fxp_sinusoid'length),
            to_signed(-5205, signed_fxp_sinusoid'length),
            to_signed(-32413, signed_fxp_sinusoid'length),
            to_signed(-4808, signed_fxp_sinusoid'length),
            to_signed(-32469, signed_fxp_sinusoid'length),
            to_signed(-4409, signed_fxp_sinusoid'length),
            to_signed(-32521, signed_fxp_sinusoid'length),
            to_signed(-4011, signed_fxp_sinusoid'length),
            to_signed(-32568, signed_fxp_sinusoid'length),
            to_signed(-3611, signed_fxp_sinusoid'length),
            to_signed(-32610, signed_fxp_sinusoid'length),
            to_signed(-3211, signed_fxp_sinusoid'length),
            to_signed(-32647, signed_fxp_sinusoid'length),
            to_signed(-2811, signed_fxp_sinusoid'length),
            to_signed(-32679, signed_fxp_sinusoid'length),
            to_signed(-2410, signed_fxp_sinusoid'length),
            to_signed(-32706, signed_fxp_sinusoid'length),
            to_signed(-2009, signed_fxp_sinusoid'length),
            to_signed(-32728, signed_fxp_sinusoid'length),
            to_signed(-1607, signed_fxp_sinusoid'length),
            to_signed(-32745, signed_fxp_sinusoid'length),
            to_signed(-1206, signed_fxp_sinusoid'length),
            to_signed(-32758, signed_fxp_sinusoid'length),
            to_signed(-804, signed_fxp_sinusoid'length),
            to_signed(-32765, signed_fxp_sinusoid'length),
            to_signed(-402, signed_fxp_sinusoid'length)
        );
end package DFTSinusoidLUT;