library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.math_real.all;

library work;
use work.DFTTypes.all;

package DFTSinusoidLUT is
    
    type sinusoid_LUT_array is   array (2*K_LENGTH-1 downto 0) of signed_fxp_sinusoid;
    
    -- format:
    -- 0: cos(-2*pi*k0/#samples)
    -- 1: sin(-2*pi*k0/#samples)
    -- 2: cos(-2*pi*k1/#samples)
    -- 3: sin(-2*pi*k1/#samples)
    -- ...

    constant K_SINUSOID_LUT   : sinusoid_LUT_array :=
        (
            -- WINDOW: 512, RESOLUTION (K-STEP): 8
            -- to_signed(32767, signed_fxp_sinusoid'length),
            -- to_signed(0, signed_fxp_sinusoid'length),
            -- to_signed(32609, signed_fxp_sinusoid'length),
            -- to_signed(-3211, signed_fxp_sinusoid'length),
            -- to_signed(32137, signed_fxp_sinusoid'length),
            -- to_signed(-6392, signed_fxp_sinusoid'length),
            -- to_signed(31356, signed_fxp_sinusoid'length),
            -- to_signed(-9511, signed_fxp_sinusoid'length),
            -- to_signed(30272, signed_fxp_sinusoid'length),
            -- to_signed(-12539, signed_fxp_sinusoid'length),
            -- to_signed(28897, signed_fxp_sinusoid'length),
            -- to_signed(-15446, signed_fxp_sinusoid'length),
            -- to_signed(27244, signed_fxp_sinusoid'length),
            -- to_signed(-18204, signed_fxp_sinusoid'length),
            -- to_signed(25329, signed_fxp_sinusoid'length),
            -- to_signed(-20787, signed_fxp_sinusoid'length),
            -- to_signed(23169, signed_fxp_sinusoid'length),
            -- to_signed(-23169, signed_fxp_sinusoid'length),
            -- to_signed(20787, signed_fxp_sinusoid'length),
            -- to_signed(-25329, signed_fxp_sinusoid'length),
            -- to_signed(18204, signed_fxp_sinusoid'length),
            -- to_signed(-27244, signed_fxp_sinusoid'length),
            -- to_signed(15446, signed_fxp_sinusoid'length),
            -- to_signed(-28897, signed_fxp_sinusoid'length),
            -- to_signed(12539, signed_fxp_sinusoid'length),
            -- to_signed(-30272, signed_fxp_sinusoid'length),
            -- to_signed(9511, signed_fxp_sinusoid'length),
            -- to_signed(-31356, signed_fxp_sinusoid'length),
            -- to_signed(6392, signed_fxp_sinusoid'length),
            -- to_signed(-32137, signed_fxp_sinusoid'length),
            -- to_signed(3211, signed_fxp_sinusoid'length),
            -- to_signed(-32609, signed_fxp_sinusoid'length),
            -- to_signed(0, signed_fxp_sinusoid'length),
            -- to_signed(-32767, signed_fxp_sinusoid'length),
            -- to_signed(-3211, signed_fxp_sinusoid'length),
            -- to_signed(-32609, signed_fxp_sinusoid'length),
            -- to_signed(-6392, signed_fxp_sinusoid'length),
            -- to_signed(-32137, signed_fxp_sinusoid'length),
            -- to_signed(-9511, signed_fxp_sinusoid'length),
            -- to_signed(-31356, signed_fxp_sinusoid'length),
            -- to_signed(-12539, signed_fxp_sinusoid'length),
            -- to_signed(-30272, signed_fxp_sinusoid'length),
            -- to_signed(-15446, signed_fxp_sinusoid'length),
            -- to_signed(-28897, signed_fxp_sinusoid'length),
            -- to_signed(-18204, signed_fxp_sinusoid'length),
            -- to_signed(-27244, signed_fxp_sinusoid'length),
            -- to_signed(-20787, signed_fxp_sinusoid'length),
            -- to_signed(-25329, signed_fxp_sinusoid'length),
            -- to_signed(-23169, signed_fxp_sinusoid'length),
            -- to_signed(-23169, signed_fxp_sinusoid'length),
            -- to_signed(-25329, signed_fxp_sinusoid'length),
            -- to_signed(-20787, signed_fxp_sinusoid'length),
            -- to_signed(-27244, signed_fxp_sinusoid'length),
            -- to_signed(-18204, signed_fxp_sinusoid'length),
            -- to_signed(-28897, signed_fxp_sinusoid'length),
            -- to_signed(-15446, signed_fxp_sinusoid'length),
            -- to_signed(-30272, signed_fxp_sinusoid'length),
            -- to_signed(-12539, signed_fxp_sinusoid'length),
            -- to_signed(-31356, signed_fxp_sinusoid'length),
            -- to_signed(-9511, signed_fxp_sinusoid'length),
            -- to_signed(-32137, signed_fxp_sinusoid'length),
            -- to_signed(-6392, signed_fxp_sinusoid'length),
            -- to_signed(-32609, signed_fxp_sinusoid'length),
            -- to_signed(-3211, signed_fxp_sinusoid'length)

            -- WINDOW: 512, RESOLUTION (K-STEP): 4
            to_signed(32767, signed_fxp_sinusoid'length),
            to_signed(0, signed_fxp_sinusoid'length),
            to_signed(32727, signed_fxp_sinusoid'length),
            to_signed(-1607, signed_fxp_sinusoid'length),
            to_signed(32609, signed_fxp_sinusoid'length),
            to_signed(-3211, signed_fxp_sinusoid'length),
            to_signed(32412, signed_fxp_sinusoid'length),
            to_signed(-4807, signed_fxp_sinusoid'length),
            to_signed(32137, signed_fxp_sinusoid'length),
            to_signed(-6392, signed_fxp_sinusoid'length),
            to_signed(31785, signed_fxp_sinusoid'length),
            to_signed(-7961, signed_fxp_sinusoid'length),
            to_signed(31356, signed_fxp_sinusoid'length),
            to_signed(-9511, signed_fxp_sinusoid'length),
            to_signed(30851, signed_fxp_sinusoid'length),
            to_signed(-11038, signed_fxp_sinusoid'length),
            to_signed(30272, signed_fxp_sinusoid'length),
            to_signed(-12539, signed_fxp_sinusoid'length),
            to_signed(29621, signed_fxp_sinusoid'length),
            to_signed(-14009, signed_fxp_sinusoid'length),
            to_signed(28897, signed_fxp_sinusoid'length),
            to_signed(-15446, signed_fxp_sinusoid'length),
            to_signed(28105, signed_fxp_sinusoid'length),
            to_signed(-16845, signed_fxp_sinusoid'length),
            to_signed(27244, signed_fxp_sinusoid'length),
            to_signed(-18204, signed_fxp_sinusoid'length),
            to_signed(26318, signed_fxp_sinusoid'length),
            to_signed(-19519, signed_fxp_sinusoid'length),
            to_signed(25329, signed_fxp_sinusoid'length),
            to_signed(-20787, signed_fxp_sinusoid'length),
            to_signed(24278, signed_fxp_sinusoid'length),
            to_signed(-22004, signed_fxp_sinusoid'length),
            to_signed(23169, signed_fxp_sinusoid'length),
            to_signed(-23169, signed_fxp_sinusoid'length),
            to_signed(22004, signed_fxp_sinusoid'length),
            to_signed(-24278, signed_fxp_sinusoid'length),
            to_signed(20787, signed_fxp_sinusoid'length),
            to_signed(-25329, signed_fxp_sinusoid'length),
            to_signed(19519, signed_fxp_sinusoid'length),
            to_signed(-26318, signed_fxp_sinusoid'length),
            to_signed(18204, signed_fxp_sinusoid'length),
            to_signed(-27244, signed_fxp_sinusoid'length),
            to_signed(16845, signed_fxp_sinusoid'length),
            to_signed(-28105, signed_fxp_sinusoid'length),
            to_signed(15446, signed_fxp_sinusoid'length),
            to_signed(-28897, signed_fxp_sinusoid'length),
            to_signed(14009, signed_fxp_sinusoid'length),
            to_signed(-29621, signed_fxp_sinusoid'length),
            to_signed(12539, signed_fxp_sinusoid'length),
            to_signed(-30272, signed_fxp_sinusoid'length),
            to_signed(11038, signed_fxp_sinusoid'length),
            to_signed(-30851, signed_fxp_sinusoid'length),
            to_signed(9511, signed_fxp_sinusoid'length),
            to_signed(-31356, signed_fxp_sinusoid'length),
            to_signed(7961, signed_fxp_sinusoid'length),
            to_signed(-31785, signed_fxp_sinusoid'length),
            to_signed(6392, signed_fxp_sinusoid'length),
            to_signed(-32137, signed_fxp_sinusoid'length),
            to_signed(4807, signed_fxp_sinusoid'length),
            to_signed(-32412, signed_fxp_sinusoid'length),
            to_signed(3211, signed_fxp_sinusoid'length),
            to_signed(-32609, signed_fxp_sinusoid'length),
            to_signed(1607, signed_fxp_sinusoid'length),
            to_signed(-32727, signed_fxp_sinusoid'length),
            to_signed(0, signed_fxp_sinusoid'length),
            to_signed(-32767, signed_fxp_sinusoid'length),
            to_signed(-1607, signed_fxp_sinusoid'length),
            to_signed(-32727, signed_fxp_sinusoid'length),
            to_signed(-3211, signed_fxp_sinusoid'length),
            to_signed(-32609, signed_fxp_sinusoid'length),
            to_signed(-4807, signed_fxp_sinusoid'length),
            to_signed(-32412, signed_fxp_sinusoid'length),
            to_signed(-6392, signed_fxp_sinusoid'length),
            to_signed(-32137, signed_fxp_sinusoid'length),
            to_signed(-7961, signed_fxp_sinusoid'length),
            to_signed(-31785, signed_fxp_sinusoid'length),
            to_signed(-9511, signed_fxp_sinusoid'length),
            to_signed(-31356, signed_fxp_sinusoid'length),
            to_signed(-11038, signed_fxp_sinusoid'length),
            to_signed(-30851, signed_fxp_sinusoid'length),
            to_signed(-12539, signed_fxp_sinusoid'length),
            to_signed(-30272, signed_fxp_sinusoid'length),
            to_signed(-14009, signed_fxp_sinusoid'length),
            to_signed(-29621, signed_fxp_sinusoid'length),
            to_signed(-15446, signed_fxp_sinusoid'length),
            to_signed(-28897, signed_fxp_sinusoid'length),
            to_signed(-16845, signed_fxp_sinusoid'length),
            to_signed(-28105, signed_fxp_sinusoid'length),
            to_signed(-18204, signed_fxp_sinusoid'length),
            to_signed(-27244, signed_fxp_sinusoid'length),
            to_signed(-19519, signed_fxp_sinusoid'length),
            to_signed(-26318, signed_fxp_sinusoid'length),
            to_signed(-20787, signed_fxp_sinusoid'length),
            to_signed(-25329, signed_fxp_sinusoid'length),
            to_signed(-22004, signed_fxp_sinusoid'length),
            to_signed(-24278, signed_fxp_sinusoid'length),
            to_signed(-23169, signed_fxp_sinusoid'length),
            to_signed(-23169, signed_fxp_sinusoid'length),
            to_signed(-24278, signed_fxp_sinusoid'length),
            to_signed(-22004, signed_fxp_sinusoid'length),
            to_signed(-25329, signed_fxp_sinusoid'length),
            to_signed(-20787, signed_fxp_sinusoid'length),
            to_signed(-26318, signed_fxp_sinusoid'length),
            to_signed(-19519, signed_fxp_sinusoid'length),
            to_signed(-27244, signed_fxp_sinusoid'length),
            to_signed(-18204, signed_fxp_sinusoid'length),
            to_signed(-28105, signed_fxp_sinusoid'length),
            to_signed(-16845, signed_fxp_sinusoid'length),
            to_signed(-28897, signed_fxp_sinusoid'length),
            to_signed(-15446, signed_fxp_sinusoid'length),
            to_signed(-29621, signed_fxp_sinusoid'length),
            to_signed(-14009, signed_fxp_sinusoid'length),
            to_signed(-30272, signed_fxp_sinusoid'length),
            to_signed(-12539, signed_fxp_sinusoid'length),
            to_signed(-30851, signed_fxp_sinusoid'length),
            to_signed(-11038, signed_fxp_sinusoid'length),
            to_signed(-31356, signed_fxp_sinusoid'length),
            to_signed(-9511, signed_fxp_sinusoid'length),
            to_signed(-31785, signed_fxp_sinusoid'length),
            to_signed(-7961, signed_fxp_sinusoid'length),
            to_signed(-32137, signed_fxp_sinusoid'length),
            to_signed(-6392, signed_fxp_sinusoid'length),
            to_signed(-32412, signed_fxp_sinusoid'length),
            to_signed(-4807, signed_fxp_sinusoid'length),
            to_signed(-32609, signed_fxp_sinusoid'length),
            to_signed(-3211, signed_fxp_sinusoid'length),
            to_signed(-32727, signed_fxp_sinusoid'length),
            to_signed(-1607, signed_fxp_sinusoid'length)

            -- WINDOW: 512, RESOLUTION (K-STEP): 1
            -- to_signed(32767, signed_fxp_sinusoid'length),
            -- to_signed(0, signed_fxp_sinusoid'length),
            -- to_signed(32764, signed_fxp_sinusoid'length),
            -- to_signed(-402, signed_fxp_sinusoid'length),
            -- to_signed(32757, signed_fxp_sinusoid'length),
            -- to_signed(-804, signed_fxp_sinusoid'length),
            -- to_signed(32744, signed_fxp_sinusoid'length),
            -- to_signed(-1206, signed_fxp_sinusoid'length),
            -- to_signed(32727, signed_fxp_sinusoid'length),
            -- to_signed(-1607, signed_fxp_sinusoid'length),
            -- to_signed(32705, signed_fxp_sinusoid'length),
            -- to_signed(-2009, signed_fxp_sinusoid'length),
            -- to_signed(32678, signed_fxp_sinusoid'length),
            -- to_signed(-2410, signed_fxp_sinusoid'length),
            -- to_signed(32646, signed_fxp_sinusoid'length),
            -- to_signed(-2811, signed_fxp_sinusoid'length),
            -- to_signed(32609, signed_fxp_sinusoid'length),
            -- to_signed(-3211, signed_fxp_sinusoid'length),
            -- to_signed(32567, signed_fxp_sinusoid'length),
            -- to_signed(-3611, signed_fxp_sinusoid'length),
            -- to_signed(32520, signed_fxp_sinusoid'length),
            -- to_signed(-4011, signed_fxp_sinusoid'length),
            -- to_signed(32468, signed_fxp_sinusoid'length),
            -- to_signed(-4409, signed_fxp_sinusoid'length),
            -- to_signed(32412, signed_fxp_sinusoid'length),
            -- to_signed(-4807, signed_fxp_sinusoid'length),
            -- to_signed(32350, signed_fxp_sinusoid'length),
            -- to_signed(-5205, signed_fxp_sinusoid'length),
            -- to_signed(32284, signed_fxp_sinusoid'length),
            -- to_signed(-5601, signed_fxp_sinusoid'length),
            -- to_signed(32213, signed_fxp_sinusoid'length),
            -- to_signed(-5997, signed_fxp_sinusoid'length),
            -- to_signed(32137, signed_fxp_sinusoid'length),
            -- to_signed(-6392, signed_fxp_sinusoid'length),
            -- to_signed(32056, signed_fxp_sinusoid'length),
            -- to_signed(-6786, signed_fxp_sinusoid'length),
            -- to_signed(31970, signed_fxp_sinusoid'length),
            -- to_signed(-7179, signed_fxp_sinusoid'length),
            -- to_signed(31880, signed_fxp_sinusoid'length),
            -- to_signed(-7571, signed_fxp_sinusoid'length),
            -- to_signed(31785, signed_fxp_sinusoid'length),
            -- to_signed(-7961, signed_fxp_sinusoid'length),
            -- to_signed(31684, signed_fxp_sinusoid'length),
            -- to_signed(-8351, signed_fxp_sinusoid'length),
            -- to_signed(31580, signed_fxp_sinusoid'length),
            -- to_signed(-8739, signed_fxp_sinusoid'length),
            -- to_signed(31470, signed_fxp_sinusoid'length),
            -- to_signed(-9126, signed_fxp_sinusoid'length),
            -- to_signed(31356, signed_fxp_sinusoid'length),
            -- to_signed(-9511, signed_fxp_sinusoid'length),
            -- to_signed(31236, signed_fxp_sinusoid'length),
            -- to_signed(-9895, signed_fxp_sinusoid'length),
            -- to_signed(31113, signed_fxp_sinusoid'length),
            -- to_signed(-10278, signed_fxp_sinusoid'length),
            -- to_signed(30984, signed_fxp_sinusoid'length),
            -- to_signed(-10659, signed_fxp_sinusoid'length),
            -- to_signed(30851, signed_fxp_sinusoid'length),
            -- to_signed(-11038, signed_fxp_sinusoid'length),
            -- to_signed(30713, signed_fxp_sinusoid'length),
            -- to_signed(-11416, signed_fxp_sinusoid'length),
            -- to_signed(30571, signed_fxp_sinusoid'length),
            -- to_signed(-11792, signed_fxp_sinusoid'length),
            -- to_signed(30424, signed_fxp_sinusoid'length),
            -- to_signed(-12166, signed_fxp_sinusoid'length),
            -- to_signed(30272, signed_fxp_sinusoid'length),
            -- to_signed(-12539, signed_fxp_sinusoid'length),
            -- to_signed(30116, signed_fxp_sinusoid'length),
            -- to_signed(-12909, signed_fxp_sinusoid'length),
            -- to_signed(29955, signed_fxp_sinusoid'length),
            -- to_signed(-13278, signed_fxp_sinusoid'length),
            -- to_signed(29790, signed_fxp_sinusoid'length),
            -- to_signed(-13645, signed_fxp_sinusoid'length),
            -- to_signed(29621, signed_fxp_sinusoid'length),
            -- to_signed(-14009, signed_fxp_sinusoid'length),
            -- to_signed(29446, signed_fxp_sinusoid'length),
            -- to_signed(-14372, signed_fxp_sinusoid'length),
            -- to_signed(29268, signed_fxp_sinusoid'length),
            -- to_signed(-14732, signed_fxp_sinusoid'length),
            -- to_signed(29085, signed_fxp_sinusoid'length),
            -- to_signed(-15090, signed_fxp_sinusoid'length),
            -- to_signed(28897, signed_fxp_sinusoid'length),
            -- to_signed(-15446, signed_fxp_sinusoid'length),
            -- to_signed(28706, signed_fxp_sinusoid'length),
            -- to_signed(-15799, signed_fxp_sinusoid'length),
            -- to_signed(28510, signed_fxp_sinusoid'length),
            -- to_signed(-16150, signed_fxp_sinusoid'length),
            -- to_signed(28309, signed_fxp_sinusoid'length),
            -- to_signed(-16499, signed_fxp_sinusoid'length),
            -- to_signed(28105, signed_fxp_sinusoid'length),
            -- to_signed(-16845, signed_fxp_sinusoid'length),
            -- to_signed(27896, signed_fxp_sinusoid'length),
            -- to_signed(-17189, signed_fxp_sinusoid'length),
            -- to_signed(27683, signed_fxp_sinusoid'length),
            -- to_signed(-17530, signed_fxp_sinusoid'length),
            -- to_signed(27466, signed_fxp_sinusoid'length),
            -- to_signed(-17868, signed_fxp_sinusoid'length),
            -- to_signed(27244, signed_fxp_sinusoid'length),
            -- to_signed(-18204, signed_fxp_sinusoid'length),
            -- to_signed(27019, signed_fxp_sinusoid'length),
            -- to_signed(-18537, signed_fxp_sinusoid'length),
            -- to_signed(26789, signed_fxp_sinusoid'length),
            -- to_signed(-18867, signed_fxp_sinusoid'length),
            -- to_signed(26556, signed_fxp_sinusoid'length),
            -- to_signed(-19194, signed_fxp_sinusoid'length),
            -- to_signed(26318, signed_fxp_sinusoid'length),
            -- to_signed(-19519, signed_fxp_sinusoid'length),
            -- to_signed(26077, signed_fxp_sinusoid'length),
            -- to_signed(-19840, signed_fxp_sinusoid'length),
            -- to_signed(25831, signed_fxp_sinusoid'length),
            -- to_signed(-20159, signed_fxp_sinusoid'length),
            -- to_signed(25582, signed_fxp_sinusoid'length),
            -- to_signed(-20474, signed_fxp_sinusoid'length),
            -- to_signed(25329, signed_fxp_sinusoid'length),
            -- to_signed(-20787, signed_fxp_sinusoid'length),
            -- to_signed(25072, signed_fxp_sinusoid'length),
            -- to_signed(-21096, signed_fxp_sinusoid'length),
            -- to_signed(24811, signed_fxp_sinusoid'length),
            -- to_signed(-21402, signed_fxp_sinusoid'length),
            -- to_signed(24546, signed_fxp_sinusoid'length),
            -- to_signed(-21705, signed_fxp_sinusoid'length),
            -- to_signed(24278, signed_fxp_sinusoid'length),
            -- to_signed(-22004, signed_fxp_sinusoid'length),
            -- to_signed(24006, signed_fxp_sinusoid'length),
            -- to_signed(-22301, signed_fxp_sinusoid'length),
            -- to_signed(23731, signed_fxp_sinusoid'length),
            -- to_signed(-22594, signed_fxp_sinusoid'length),
            -- to_signed(23452, signed_fxp_sinusoid'length),
            -- to_signed(-22883, signed_fxp_sinusoid'length),
            -- to_signed(23169, signed_fxp_sinusoid'length),
            -- to_signed(-23169, signed_fxp_sinusoid'length),
            -- to_signed(22883, signed_fxp_sinusoid'length),
            -- to_signed(-23452, signed_fxp_sinusoid'length),
            -- to_signed(22594, signed_fxp_sinusoid'length),
            -- to_signed(-23731, signed_fxp_sinusoid'length),
            -- to_signed(22301, signed_fxp_sinusoid'length),
            -- to_signed(-24006, signed_fxp_sinusoid'length),
            -- to_signed(22004, signed_fxp_sinusoid'length),
            -- to_signed(-24278, signed_fxp_sinusoid'length),
            -- to_signed(21705, signed_fxp_sinusoid'length),
            -- to_signed(-24546, signed_fxp_sinusoid'length),
            -- to_signed(21402, signed_fxp_sinusoid'length),
            -- to_signed(-24811, signed_fxp_sinusoid'length),
            -- to_signed(21096, signed_fxp_sinusoid'length),
            -- to_signed(-25072, signed_fxp_sinusoid'length),
            -- to_signed(20787, signed_fxp_sinusoid'length),
            -- to_signed(-25329, signed_fxp_sinusoid'length),
            -- to_signed(20474, signed_fxp_sinusoid'length),
            -- to_signed(-25582, signed_fxp_sinusoid'length),
            -- to_signed(20159, signed_fxp_sinusoid'length),
            -- to_signed(-25831, signed_fxp_sinusoid'length),
            -- to_signed(19840, signed_fxp_sinusoid'length),
            -- to_signed(-26077, signed_fxp_sinusoid'length),
            -- to_signed(19519, signed_fxp_sinusoid'length),
            -- to_signed(-26318, signed_fxp_sinusoid'length),
            -- to_signed(19194, signed_fxp_sinusoid'length),
            -- to_signed(-26556, signed_fxp_sinusoid'length),
            -- to_signed(18867, signed_fxp_sinusoid'length),
            -- to_signed(-26789, signed_fxp_sinusoid'length),
            -- to_signed(18537, signed_fxp_sinusoid'length),
            -- to_signed(-27019, signed_fxp_sinusoid'length),
            -- to_signed(18204, signed_fxp_sinusoid'length),
            -- to_signed(-27244, signed_fxp_sinusoid'length),
            -- to_signed(17868, signed_fxp_sinusoid'length),
            -- to_signed(-27466, signed_fxp_sinusoid'length),
            -- to_signed(17530, signed_fxp_sinusoid'length),
            -- to_signed(-27683, signed_fxp_sinusoid'length),
            -- to_signed(17189, signed_fxp_sinusoid'length),
            -- to_signed(-27896, signed_fxp_sinusoid'length),
            -- to_signed(16845, signed_fxp_sinusoid'length),
            -- to_signed(-28105, signed_fxp_sinusoid'length),
            -- to_signed(16499, signed_fxp_sinusoid'length),
            -- to_signed(-28309, signed_fxp_sinusoid'length),
            -- to_signed(16150, signed_fxp_sinusoid'length),
            -- to_signed(-28510, signed_fxp_sinusoid'length),
            -- to_signed(15799, signed_fxp_sinusoid'length),
            -- to_signed(-28706, signed_fxp_sinusoid'length),
            -- to_signed(15446, signed_fxp_sinusoid'length),
            -- to_signed(-28897, signed_fxp_sinusoid'length),
            -- to_signed(15090, signed_fxp_sinusoid'length),
            -- to_signed(-29085, signed_fxp_sinusoid'length),
            -- to_signed(14732, signed_fxp_sinusoid'length),
            -- to_signed(-29268, signed_fxp_sinusoid'length),
            -- to_signed(14372, signed_fxp_sinusoid'length),
            -- to_signed(-29446, signed_fxp_sinusoid'length),
            -- to_signed(14009, signed_fxp_sinusoid'length),
            -- to_signed(-29621, signed_fxp_sinusoid'length),
            -- to_signed(13645, signed_fxp_sinusoid'length),
            -- to_signed(-29790, signed_fxp_sinusoid'length),
            -- to_signed(13278, signed_fxp_sinusoid'length),
            -- to_signed(-29955, signed_fxp_sinusoid'length),
            -- to_signed(12909, signed_fxp_sinusoid'length),
            -- to_signed(-30116, signed_fxp_sinusoid'length),
            -- to_signed(12539, signed_fxp_sinusoid'length),
            -- to_signed(-30272, signed_fxp_sinusoid'length),
            -- to_signed(12166, signed_fxp_sinusoid'length),
            -- to_signed(-30424, signed_fxp_sinusoid'length),
            -- to_signed(11792, signed_fxp_sinusoid'length),
            -- to_signed(-30571, signed_fxp_sinusoid'length),
            -- to_signed(11416, signed_fxp_sinusoid'length),
            -- to_signed(-30713, signed_fxp_sinusoid'length),
            -- to_signed(11038, signed_fxp_sinusoid'length),
            -- to_signed(-30851, signed_fxp_sinusoid'length),
            -- to_signed(10659, signed_fxp_sinusoid'length),
            -- to_signed(-30984, signed_fxp_sinusoid'length),
            -- to_signed(10278, signed_fxp_sinusoid'length),
            -- to_signed(-31113, signed_fxp_sinusoid'length),
            -- to_signed(9895, signed_fxp_sinusoid'length),
            -- to_signed(-31236, signed_fxp_sinusoid'length),
            -- to_signed(9511, signed_fxp_sinusoid'length),
            -- to_signed(-31356, signed_fxp_sinusoid'length),
            -- to_signed(9126, signed_fxp_sinusoid'length),
            -- to_signed(-31470, signed_fxp_sinusoid'length),
            -- to_signed(8739, signed_fxp_sinusoid'length),
            -- to_signed(-31580, signed_fxp_sinusoid'length),
            -- to_signed(8351, signed_fxp_sinusoid'length),
            -- to_signed(-31684, signed_fxp_sinusoid'length),
            -- to_signed(7961, signed_fxp_sinusoid'length),
            -- to_signed(-31785, signed_fxp_sinusoid'length),
            -- to_signed(7571, signed_fxp_sinusoid'length),
            -- to_signed(-31880, signed_fxp_sinusoid'length),
            -- to_signed(7179, signed_fxp_sinusoid'length),
            -- to_signed(-31970, signed_fxp_sinusoid'length),
            -- to_signed(6786, signed_fxp_sinusoid'length),
            -- to_signed(-32056, signed_fxp_sinusoid'length),
            -- to_signed(6392, signed_fxp_sinusoid'length),
            -- to_signed(-32137, signed_fxp_sinusoid'length),
            -- to_signed(5997, signed_fxp_sinusoid'length),
            -- to_signed(-32213, signed_fxp_sinusoid'length),
            -- to_signed(5601, signed_fxp_sinusoid'length),
            -- to_signed(-32284, signed_fxp_sinusoid'length),
            -- to_signed(5205, signed_fxp_sinusoid'length),
            -- to_signed(-32350, signed_fxp_sinusoid'length),
            -- to_signed(4807, signed_fxp_sinusoid'length),
            -- to_signed(-32412, signed_fxp_sinusoid'length),
            -- to_signed(4409, signed_fxp_sinusoid'length),
            -- to_signed(-32468, signed_fxp_sinusoid'length),
            -- to_signed(4011, signed_fxp_sinusoid'length),
            -- to_signed(-32520, signed_fxp_sinusoid'length),
            -- to_signed(3611, signed_fxp_sinusoid'length),
            -- to_signed(-32567, signed_fxp_sinusoid'length),
            -- to_signed(3211, signed_fxp_sinusoid'length),
            -- to_signed(-32609, signed_fxp_sinusoid'length),
            -- to_signed(2811, signed_fxp_sinusoid'length),
            -- to_signed(-32646, signed_fxp_sinusoid'length),
            -- to_signed(2410, signed_fxp_sinusoid'length),
            -- to_signed(-32678, signed_fxp_sinusoid'length),
            -- to_signed(2009, signed_fxp_sinusoid'length),
            -- to_signed(-32705, signed_fxp_sinusoid'length),
            -- to_signed(1607, signed_fxp_sinusoid'length),
            -- to_signed(-32727, signed_fxp_sinusoid'length),
            -- to_signed(1206, signed_fxp_sinusoid'length),
            -- to_signed(-32744, signed_fxp_sinusoid'length),
            -- to_signed(804, signed_fxp_sinusoid'length),
            -- to_signed(-32757, signed_fxp_sinusoid'length),
            -- to_signed(402, signed_fxp_sinusoid'length),
            -- to_signed(-32764, signed_fxp_sinusoid'length),
            -- to_signed(0, signed_fxp_sinusoid'length),
            -- to_signed(-32767, signed_fxp_sinusoid'length),
            -- to_signed(-402, signed_fxp_sinusoid'length),
            -- to_signed(-32764, signed_fxp_sinusoid'length),
            -- to_signed(-804, signed_fxp_sinusoid'length),
            -- to_signed(-32757, signed_fxp_sinusoid'length),
            -- to_signed(-1206, signed_fxp_sinusoid'length),
            -- to_signed(-32744, signed_fxp_sinusoid'length),
            -- to_signed(-1607, signed_fxp_sinusoid'length),
            -- to_signed(-32727, signed_fxp_sinusoid'length),
            -- to_signed(-2009, signed_fxp_sinusoid'length),
            -- to_signed(-32705, signed_fxp_sinusoid'length),
            -- to_signed(-2410, signed_fxp_sinusoid'length),
            -- to_signed(-32678, signed_fxp_sinusoid'length),
            -- to_signed(-2811, signed_fxp_sinusoid'length),
            -- to_signed(-32646, signed_fxp_sinusoid'length),
            -- to_signed(-3211, signed_fxp_sinusoid'length),
            -- to_signed(-32609, signed_fxp_sinusoid'length),
            -- to_signed(-3611, signed_fxp_sinusoid'length),
            -- to_signed(-32567, signed_fxp_sinusoid'length),
            -- to_signed(-4011, signed_fxp_sinusoid'length),
            -- to_signed(-32520, signed_fxp_sinusoid'length),
            -- to_signed(-4409, signed_fxp_sinusoid'length),
            -- to_signed(-32468, signed_fxp_sinusoid'length),
            -- to_signed(-4807, signed_fxp_sinusoid'length),
            -- to_signed(-32412, signed_fxp_sinusoid'length),
            -- to_signed(-5205, signed_fxp_sinusoid'length),
            -- to_signed(-32350, signed_fxp_sinusoid'length),
            -- to_signed(-5601, signed_fxp_sinusoid'length),
            -- to_signed(-32284, signed_fxp_sinusoid'length),
            -- to_signed(-5997, signed_fxp_sinusoid'length),
            -- to_signed(-32213, signed_fxp_sinusoid'length),
            -- to_signed(-6392, signed_fxp_sinusoid'length),
            -- to_signed(-32137, signed_fxp_sinusoid'length),
            -- to_signed(-6786, signed_fxp_sinusoid'length),
            -- to_signed(-32056, signed_fxp_sinusoid'length),
            -- to_signed(-7179, signed_fxp_sinusoid'length),
            -- to_signed(-31970, signed_fxp_sinusoid'length),
            -- to_signed(-7571, signed_fxp_sinusoid'length),
            -- to_signed(-31880, signed_fxp_sinusoid'length),
            -- to_signed(-7961, signed_fxp_sinusoid'length),
            -- to_signed(-31785, signed_fxp_sinusoid'length),
            -- to_signed(-8351, signed_fxp_sinusoid'length),
            -- to_signed(-31684, signed_fxp_sinusoid'length),
            -- to_signed(-8739, signed_fxp_sinusoid'length),
            -- to_signed(-31580, signed_fxp_sinusoid'length),
            -- to_signed(-9126, signed_fxp_sinusoid'length),
            -- to_signed(-31470, signed_fxp_sinusoid'length),
            -- to_signed(-9511, signed_fxp_sinusoid'length),
            -- to_signed(-31356, signed_fxp_sinusoid'length),
            -- to_signed(-9895, signed_fxp_sinusoid'length),
            -- to_signed(-31236, signed_fxp_sinusoid'length),
            -- to_signed(-10278, signed_fxp_sinusoid'length),
            -- to_signed(-31113, signed_fxp_sinusoid'length),
            -- to_signed(-10659, signed_fxp_sinusoid'length),
            -- to_signed(-30984, signed_fxp_sinusoid'length),
            -- to_signed(-11038, signed_fxp_sinusoid'length),
            -- to_signed(-30851, signed_fxp_sinusoid'length),
            -- to_signed(-11416, signed_fxp_sinusoid'length),
            -- to_signed(-30713, signed_fxp_sinusoid'length),
            -- to_signed(-11792, signed_fxp_sinusoid'length),
            -- to_signed(-30571, signed_fxp_sinusoid'length),
            -- to_signed(-12166, signed_fxp_sinusoid'length),
            -- to_signed(-30424, signed_fxp_sinusoid'length),
            -- to_signed(-12539, signed_fxp_sinusoid'length),
            -- to_signed(-30272, signed_fxp_sinusoid'length),
            -- to_signed(-12909, signed_fxp_sinusoid'length),
            -- to_signed(-30116, signed_fxp_sinusoid'length),
            -- to_signed(-13278, signed_fxp_sinusoid'length),
            -- to_signed(-29955, signed_fxp_sinusoid'length),
            -- to_signed(-13645, signed_fxp_sinusoid'length),
            -- to_signed(-29790, signed_fxp_sinusoid'length),
            -- to_signed(-14009, signed_fxp_sinusoid'length),
            -- to_signed(-29621, signed_fxp_sinusoid'length),
            -- to_signed(-14372, signed_fxp_sinusoid'length),
            -- to_signed(-29446, signed_fxp_sinusoid'length),
            -- to_signed(-14732, signed_fxp_sinusoid'length),
            -- to_signed(-29268, signed_fxp_sinusoid'length),
            -- to_signed(-15090, signed_fxp_sinusoid'length),
            -- to_signed(-29085, signed_fxp_sinusoid'length),
            -- to_signed(-15446, signed_fxp_sinusoid'length),
            -- to_signed(-28897, signed_fxp_sinusoid'length),
            -- to_signed(-15799, signed_fxp_sinusoid'length),
            -- to_signed(-28706, signed_fxp_sinusoid'length),
            -- to_signed(-16150, signed_fxp_sinusoid'length),
            -- to_signed(-28510, signed_fxp_sinusoid'length),
            -- to_signed(-16499, signed_fxp_sinusoid'length),
            -- to_signed(-28309, signed_fxp_sinusoid'length),
            -- to_signed(-16845, signed_fxp_sinusoid'length),
            -- to_signed(-28105, signed_fxp_sinusoid'length),
            -- to_signed(-17189, signed_fxp_sinusoid'length),
            -- to_signed(-27896, signed_fxp_sinusoid'length),
            -- to_signed(-17530, signed_fxp_sinusoid'length),
            -- to_signed(-27683, signed_fxp_sinusoid'length),
            -- to_signed(-17868, signed_fxp_sinusoid'length),
            -- to_signed(-27466, signed_fxp_sinusoid'length),
            -- to_signed(-18204, signed_fxp_sinusoid'length),
            -- to_signed(-27244, signed_fxp_sinusoid'length),
            -- to_signed(-18537, signed_fxp_sinusoid'length),
            -- to_signed(-27019, signed_fxp_sinusoid'length),
            -- to_signed(-18867, signed_fxp_sinusoid'length),
            -- to_signed(-26789, signed_fxp_sinusoid'length),
            -- to_signed(-19194, signed_fxp_sinusoid'length),
            -- to_signed(-26556, signed_fxp_sinusoid'length),
            -- to_signed(-19519, signed_fxp_sinusoid'length),
            -- to_signed(-26318, signed_fxp_sinusoid'length),
            -- to_signed(-19840, signed_fxp_sinusoid'length),
            -- to_signed(-26077, signed_fxp_sinusoid'length),
            -- to_signed(-20159, signed_fxp_sinusoid'length),
            -- to_signed(-25831, signed_fxp_sinusoid'length),
            -- to_signed(-20474, signed_fxp_sinusoid'length),
            -- to_signed(-25582, signed_fxp_sinusoid'length),
            -- to_signed(-20787, signed_fxp_sinusoid'length),
            -- to_signed(-25329, signed_fxp_sinusoid'length),
            -- to_signed(-21096, signed_fxp_sinusoid'length),
            -- to_signed(-25072, signed_fxp_sinusoid'length),
            -- to_signed(-21402, signed_fxp_sinusoid'length),
            -- to_signed(-24811, signed_fxp_sinusoid'length),
            -- to_signed(-21705, signed_fxp_sinusoid'length),
            -- to_signed(-24546, signed_fxp_sinusoid'length),
            -- to_signed(-22004, signed_fxp_sinusoid'length),
            -- to_signed(-24278, signed_fxp_sinusoid'length),
            -- to_signed(-22301, signed_fxp_sinusoid'length),
            -- to_signed(-24006, signed_fxp_sinusoid'length),
            -- to_signed(-22594, signed_fxp_sinusoid'length),
            -- to_signed(-23731, signed_fxp_sinusoid'length),
            -- to_signed(-22883, signed_fxp_sinusoid'length),
            -- to_signed(-23452, signed_fxp_sinusoid'length),
            -- to_signed(-23169, signed_fxp_sinusoid'length),
            -- to_signed(-23169, signed_fxp_sinusoid'length),
            -- to_signed(-23452, signed_fxp_sinusoid'length),
            -- to_signed(-22883, signed_fxp_sinusoid'length),
            -- to_signed(-23731, signed_fxp_sinusoid'length),
            -- to_signed(-22594, signed_fxp_sinusoid'length),
            -- to_signed(-24006, signed_fxp_sinusoid'length),
            -- to_signed(-22301, signed_fxp_sinusoid'length),
            -- to_signed(-24278, signed_fxp_sinusoid'length),
            -- to_signed(-22004, signed_fxp_sinusoid'length),
            -- to_signed(-24546, signed_fxp_sinusoid'length),
            -- to_signed(-21705, signed_fxp_sinusoid'length),
            -- to_signed(-24811, signed_fxp_sinusoid'length),
            -- to_signed(-21402, signed_fxp_sinusoid'length),
            -- to_signed(-25072, signed_fxp_sinusoid'length),
            -- to_signed(-21096, signed_fxp_sinusoid'length),
            -- to_signed(-25329, signed_fxp_sinusoid'length),
            -- to_signed(-20787, signed_fxp_sinusoid'length),
            -- to_signed(-25582, signed_fxp_sinusoid'length),
            -- to_signed(-20474, signed_fxp_sinusoid'length),
            -- to_signed(-25831, signed_fxp_sinusoid'length),
            -- to_signed(-20159, signed_fxp_sinusoid'length),
            -- to_signed(-26077, signed_fxp_sinusoid'length),
            -- to_signed(-19840, signed_fxp_sinusoid'length),
            -- to_signed(-26318, signed_fxp_sinusoid'length),
            -- to_signed(-19519, signed_fxp_sinusoid'length),
            -- to_signed(-26556, signed_fxp_sinusoid'length),
            -- to_signed(-19194, signed_fxp_sinusoid'length),
            -- to_signed(-26789, signed_fxp_sinusoid'length),
            -- to_signed(-18867, signed_fxp_sinusoid'length),
            -- to_signed(-27019, signed_fxp_sinusoid'length),
            -- to_signed(-18537, signed_fxp_sinusoid'length),
            -- to_signed(-27244, signed_fxp_sinusoid'length),
            -- to_signed(-18204, signed_fxp_sinusoid'length),
            -- to_signed(-27466, signed_fxp_sinusoid'length),
            -- to_signed(-17868, signed_fxp_sinusoid'length),
            -- to_signed(-27683, signed_fxp_sinusoid'length),
            -- to_signed(-17530, signed_fxp_sinusoid'length),
            -- to_signed(-27896, signed_fxp_sinusoid'length),
            -- to_signed(-17189, signed_fxp_sinusoid'length),
            -- to_signed(-28105, signed_fxp_sinusoid'length),
            -- to_signed(-16845, signed_fxp_sinusoid'length),
            -- to_signed(-28309, signed_fxp_sinusoid'length),
            -- to_signed(-16499, signed_fxp_sinusoid'length),
            -- to_signed(-28510, signed_fxp_sinusoid'length),
            -- to_signed(-16150, signed_fxp_sinusoid'length),
            -- to_signed(-28706, signed_fxp_sinusoid'length),
            -- to_signed(-15799, signed_fxp_sinusoid'length),
            -- to_signed(-28897, signed_fxp_sinusoid'length),
            -- to_signed(-15446, signed_fxp_sinusoid'length),
            -- to_signed(-29085, signed_fxp_sinusoid'length),
            -- to_signed(-15090, signed_fxp_sinusoid'length),
            -- to_signed(-29268, signed_fxp_sinusoid'length),
            -- to_signed(-14732, signed_fxp_sinusoid'length),
            -- to_signed(-29446, signed_fxp_sinusoid'length),
            -- to_signed(-14372, signed_fxp_sinusoid'length),
            -- to_signed(-29621, signed_fxp_sinusoid'length),
            -- to_signed(-14009, signed_fxp_sinusoid'length),
            -- to_signed(-29790, signed_fxp_sinusoid'length),
            -- to_signed(-13645, signed_fxp_sinusoid'length),
            -- to_signed(-29955, signed_fxp_sinusoid'length),
            -- to_signed(-13278, signed_fxp_sinusoid'length),
            -- to_signed(-30116, signed_fxp_sinusoid'length),
            -- to_signed(-12909, signed_fxp_sinusoid'length),
            -- to_signed(-30272, signed_fxp_sinusoid'length),
            -- to_signed(-12539, signed_fxp_sinusoid'length),
            -- to_signed(-30424, signed_fxp_sinusoid'length),
            -- to_signed(-12166, signed_fxp_sinusoid'length),
            -- to_signed(-30571, signed_fxp_sinusoid'length),
            -- to_signed(-11792, signed_fxp_sinusoid'length),
            -- to_signed(-30713, signed_fxp_sinusoid'length),
            -- to_signed(-11416, signed_fxp_sinusoid'length),
            -- to_signed(-30851, signed_fxp_sinusoid'length),
            -- to_signed(-11038, signed_fxp_sinusoid'length),
            -- to_signed(-30984, signed_fxp_sinusoid'length),
            -- to_signed(-10659, signed_fxp_sinusoid'length),
            -- to_signed(-31113, signed_fxp_sinusoid'length),
            -- to_signed(-10278, signed_fxp_sinusoid'length),
            -- to_signed(-31236, signed_fxp_sinusoid'length),
            -- to_signed(-9895, signed_fxp_sinusoid'length),
            -- to_signed(-31356, signed_fxp_sinusoid'length),
            -- to_signed(-9511, signed_fxp_sinusoid'length),
            -- to_signed(-31470, signed_fxp_sinusoid'length),
            -- to_signed(-9126, signed_fxp_sinusoid'length),
            -- to_signed(-31580, signed_fxp_sinusoid'length),
            -- to_signed(-8739, signed_fxp_sinusoid'length),
            -- to_signed(-31684, signed_fxp_sinusoid'length),
            -- to_signed(-8351, signed_fxp_sinusoid'length),
            -- to_signed(-31785, signed_fxp_sinusoid'length),
            -- to_signed(-7961, signed_fxp_sinusoid'length),
            -- to_signed(-31880, signed_fxp_sinusoid'length),
            -- to_signed(-7571, signed_fxp_sinusoid'length),
            -- to_signed(-31970, signed_fxp_sinusoid'length),
            -- to_signed(-7179, signed_fxp_sinusoid'length),
            -- to_signed(-32056, signed_fxp_sinusoid'length),
            -- to_signed(-6786, signed_fxp_sinusoid'length),
            -- to_signed(-32137, signed_fxp_sinusoid'length),
            -- to_signed(-6392, signed_fxp_sinusoid'length),
            -- to_signed(-32213, signed_fxp_sinusoid'length),
            -- to_signed(-5997, signed_fxp_sinusoid'length),
            -- to_signed(-32284, signed_fxp_sinusoid'length),
            -- to_signed(-5601, signed_fxp_sinusoid'length),
            -- to_signed(-32350, signed_fxp_sinusoid'length),
            -- to_signed(-5205, signed_fxp_sinusoid'length),
            -- to_signed(-32412, signed_fxp_sinusoid'length),
            -- to_signed(-4807, signed_fxp_sinusoid'length),
            -- to_signed(-32468, signed_fxp_sinusoid'length),
            -- to_signed(-4409, signed_fxp_sinusoid'length),
            -- to_signed(-32520, signed_fxp_sinusoid'length),
            -- to_signed(-4011, signed_fxp_sinusoid'length),
            -- to_signed(-32567, signed_fxp_sinusoid'length),
            -- to_signed(-3611, signed_fxp_sinusoid'length),
            -- to_signed(-32609, signed_fxp_sinusoid'length),
            -- to_signed(-3211, signed_fxp_sinusoid'length),
            -- to_signed(-32646, signed_fxp_sinusoid'length),
            -- to_signed(-2811, signed_fxp_sinusoid'length),
            -- to_signed(-32678, signed_fxp_sinusoid'length),
            -- to_signed(-2410, signed_fxp_sinusoid'length),
            -- to_signed(-32705, signed_fxp_sinusoid'length),
            -- to_signed(-2009, signed_fxp_sinusoid'length),
            -- to_signed(-32727, signed_fxp_sinusoid'length),
            -- to_signed(-1607, signed_fxp_sinusoid'length),
            -- to_signed(-32744, signed_fxp_sinusoid'length),
            -- to_signed(-1206, signed_fxp_sinusoid'length),
            -- to_signed(-32757, signed_fxp_sinusoid'length),
            -- to_signed(-804, signed_fxp_sinusoid'length),
            -- to_signed(-32764, signed_fxp_sinusoid'length),
            -- to_signed(-402, signed_fxp_sinusoid'length)
        );
end package DFTSinusoidLUT;